library verilog;
use verilog.vl_types.all;
entity ALU is
end ALU;
