library verilog;
use verilog.vl_types.all;
entity tb_L1_D_controller is
end tb_L1_D_controller;
