`timescale 1ns/100ps

module tb_ALU;
ALU u_ALU ();

endmodule